//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO
// Engineer:  Edgar Barba & Jorge Velazquez
// Module: RegisterFile
// Description: 
// Set of 32 Register for multiple purposes with selector and write control.
// 
//////////////////////////////////////////////////////////////////////////////////
module RegisterFile #(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=5)(
  input clk,
  input rst,
  input we3,
  input [(ADDR_WIDTH-1):0] A1,
  input [(ADDR_WIDTH-1):0] A2,
  input [(ADDR_WIDTH-1):0] A3,
  input [(DATA_WIDTH-1):0] wd3,
  output [(DATA_WIDTH-1):0] rd1,
  output [(DATA_WIDTH-1):0] rd2
);

wire [DATA_WIDTH-1:0] Q [2**ADDR_WIDTH-1:0]; //Declaration for all the output wires of each Register.
wire en [DATA_WIDTH-1:0]; //Declaration for all enable wires of each Register.

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Write control Module.
WriteControl WC_32_regs (
.sel(A3),
.en(we3),
.out0(en[0]),
.out1(en[1]),
.out2(en[2]),
.out3(en[3]),
.out4(en[4]),
.out5(en[5]),
.out6(en[6]),
.out7(en[7]),
.out8(en[8]),
.out9(en[9]),
.out10(en[10]),
.out11(en[11]),
.out12(en[12]),
.out13(en[13]),
.out14(en[14]),
.out15(en[15]),
.out16(en[16]),
.out17(en[17]),
.out18(en[18]),
.out19(en[19]),
.out20(en[20]),
.out21(en[21]),
.out22(en[22]),
.out23(en[23]),
.out24(en[24]),
.out25(en[25]),
.out26(en[26]),
.out27(en[27]),
.out28(en[28]),
.out29(en[29]),
.out30(en[30]),
.out31(en[31])
);
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Registers declaration.
Registers Regs (
 .D(wd3),
 .clk(clk),
 .rst(rst),
 .en0(1'b0),
 .en1(en[1]),
 .en2(en[2]),
 .en3(en[3]),
 .en4(en[4]),
 .en5(en[5]),
 .en6(en[6]),
 .en7(en[7]),
 .en8(en[8]),
 .en9(en[9]),
 .en10(en[10]),
 .en11(en[11]),
 .en12(en[12]),
 .en13(en[13]),
 .en14(en[14]),
 .en15(en[15]),
 .en16(en[16]),
 .en17(en[17]),
 .en18(en[18]),
 .en19(en[19]),
 .en20(en[20]),
 .en21(en[21]),
 .en22(en[22]),
 .en23(en[23]),
 .en24(en[24]),
 .en25(en[25]),
 .en26(en[26]),
 .en27(en[27]),
 .en28(en[28]),
 .en29(en[29]),
 .en30(en[30]),
 .en31(en[31]),
 .Q0(Q[0]),
 .Q1(Q[1]),
 .Q2(Q[2]),
 .Q3(Q[3]),
 .Q4(Q[4]),
 .Q5(Q[5]),
 .Q6(Q[6]),
 .Q7(Q[7]),
 .Q8(Q[8]),
 .Q9(Q[9]),
 .Q10(Q[10]),
 .Q11(Q[11]),
 .Q12(Q[12]),
 .Q13(Q[13]),
 .Q14(Q[14]),
 .Q15(Q[15]),
 .Q16(Q[16]),
 .Q17(Q[17]),
 .Q18(Q[18]),
 .Q19(Q[19]),
 .Q20(Q[20]),
 .Q21(Q[21]),
 .Q22(Q[22]),
 .Q23(Q[23]),
 .Q24(Q[24]),
 .Q25(Q[25]),
 .Q26(Q[26]),
 .Q27(Q[27]),
 .Q28(Q[28]),
 .Q29(Q[29]),
 .Q30(Q[30]),
 .Q31(Q[31])
);
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//32 to 1 Output MUX for RD1 selection.
MUX32input rd1Out(
  .sel(A1),
  .Q0(Q[0]),
  .Q1(Q[1]),
  .Q2(Q[2]),
  .Q3(Q[3]),
  .Q4(Q[4]),
  .Q5(Q[5]),
  .Q6(Q[6]),
  .Q7(Q[7]),
  .Q8(Q[8]),
  .Q9(Q[9]),
  .Q10(Q[10]),
  .Q11(Q[11]),
  .Q12(Q[12]),
  .Q13(Q[13]),
  .Q14(Q[14]),
  .Q15(Q[15]),
  .Q16(Q[16]),
  .Q17(Q[17]),
  .Q18(Q[18]),
  .Q19(Q[19]),
  .Q20(Q[20]),
  .Q21(Q[21]),
  .Q22(Q[22]),
  .Q23(Q[23]),
  .Q24(Q[24]),
  .Q25(Q[25]),
  .Q26(Q[26]),
  .Q27(Q[27]),
  .Q28(Q[28]),
  .Q29(Q[29]),
  .Q30(Q[30]),
  .Q31(Q[31]),
  .data(rd1)
);
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//32 to 1 Output MUX for RD2 selection.
MUX32input rd2Out(
  .sel(A2),
  .Q0(Q[0]),
  .Q1(Q[1]),
  .Q2(Q[2]),
  .Q3(Q[3]),
  .Q4(Q[4]),
  .Q5(Q[5]),
  .Q6(Q[6]),
  .Q7(Q[7]),
  .Q8(Q[8]),
  .Q9(Q[9]),
  .Q10(Q[10]),
  .Q11(Q[11]),
  .Q12(Q[12]),
  .Q13(Q[13]),
  .Q14(Q[14]),
  .Q15(Q[15]),
  .Q16(Q[16]),
  .Q17(Q[17]),
  .Q18(Q[18]),
  .Q19(Q[19]),
  .Q20(Q[20]),
  .Q21(Q[21]),
  .Q22(Q[22]),
  .Q23(Q[23]),
  .Q24(Q[24]),
  .Q25(Q[25]),
  .Q26(Q[26]),
  .Q27(Q[27]),
  .Q28(Q[28]),
  .Q29(Q[29]),
  .Q30(Q[30]),
  .Q31(Q[31]),
  .data(rd2)
);

endmodule
